module selector (input 