module manual_control_rele(clk);
input clk;


always @(posedge clk) begin
	
	
	
end

endmodule